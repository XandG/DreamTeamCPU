LIBRARY ieee;
USE ieee.std_logic_1164.all; 

ENTITY bus_phase1 IS 
	PORT(
	r0, r1, r2, r3, r4, r5, r6, r7, r8, r9, r10, r11, r12, r13, r14,
	r15, hi, lo, z_hi, z_lo, pc, mdr, inport, c_sign_extended   : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	input: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	output : OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
END bus_phase1;

ARCHITECTURE description OF bus_phase1 IS 

COMPONENT encoder32to5 
PORT(
    input: IN STD_LOGIC_VECTOR(31 DOWNTO 0);	--generated by control
    sel : OUT STD_LOGIC_VECTOR(4 DOWNTO 0) -- internal selet
	);
END COMPONENT;

COMPONENT bus_mux_24to5
 PORT(
    r0, r1, r2, r3, r4, r5, r6, r7, r8, r9, r10, r11, r12, r13, r14, r15, hi, lo, z_hi, z_lo, pc, mdr, inport, c_sign_extended   : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	 s_in : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
	 output : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END COMPONENT;

COMPONENT reg32bit
 PORT(
    d   : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    ld  : IN STD_LOGIC; -- load/enable.
    rst_n : IN STD_LOGIC; -- async. clear.
    clk : IN STD_LOGIC; -- clock.
    q   : OUT STD_LOGIC_VECTOR(31 DOWNTO 0) -- output
);
END COMPONENT;
COMPONENT MDR_unit
	PORT(
		read_sel :  IN  STD_LOGIC;
		ld :  IN  STD_LOGIC;
		rst_n :  IN  STD_LOGIC;
		clk :  IN  STD_LOGIC;
		BusMuxOut :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		MDataIn :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		Bus_Mux_In :  OUT  STD_LOGIC_VECTOR(31 DOWNTO 0));
END COMPONENT;




SIGNAL in_sig: STD_LOGIC_VECTOR(31 DOWNTO 0); --generated by control
SIGNAL out_sig: STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL r0_s, r1_s, r2_s, r3_s, r4_s, r5_s, r6_s, r7_s, r8_s, r9_s, r10_s, r11_s, 
		 r12_s, r13_s, r14_s, r15_s, hi_s, lo_s, z_hi_s, z_lo_s, pc_s, mdr_s, inport_s,
		 c_sign_extended_s   : STD_LOGIC_VECTOR(31 DOWNTO 0);
		

SIGNAL sel: STD_LOGIC_VECTOR(4 DOWNTO 0);--Internal signal
--register signals
SIGNAL q00_s, q01_s, q02_s, q03_s, q04_s, q05_s, q06_s, q07_s, q08_s, 
		 q09_s, q10_s, q11_s, q12_s, q13_s, q14_s, q15_s, q_hi_s, q_lo_s,
		 q_z_hi_s, q_z_lo_s, q_pc_s, q_mdr_s, q_inport_s, q_c_sign_extended_s	
		 :STD_LOGIC_VECTOR(31 DOWNTO 0);

SIGNAL ld00_s, ld01_s, ld02_s, ld03_s, ld04_s, ld05_s, ld06_s, ld07_s, ld08_s, 
		 ld09_s, ld10_s, ld11_s, ld12_s, ld13_s, ld14_s, ld15_s, ld_hi_s, ld_lo_s,
		 ld_z_hi_s, ld_z_lo_s, ld_pc_s, ld_mdr_s, ld_inport_s, ld_c_sign_extended_s	
		 :STD_LOGIC;
		 

--control generated global signals
SIGNAL clk_s: STD_LOGIC;
SIGNAL rst_n_s: STD_LOGIC;
--control generated MDR signals
SIGNAL Mdatain_s: STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL read_sel_s: STD_LOGIC;



BEGIN
encoder: encoder32to5
	PORT MAP(
	input=>in_sig, --generated by control 
	sel=>sel);
	
mux:bus_mux_24to5
	PORT MAP(
	r0=>q00_s,--inputs from register outputs
	r1=>q01_s,
	r2=>q02_s,
	r3=>q03_s,
	r4=>q04_s,
	r5=>q05_s,
	r6=>q06_s,
	r7=>q07_s,
	r8=>q08_s,
	r9=>q09_s,
	r10=>q10_s,
	r11=>q11_s,
	r12=>q12_s,
	r13=>q13_s,
	r14=>q14_s,
	r15=>q15_s,
	hi=>q_hi_s,
	lo=>q_lo_s,
	z_hi=>q_z_hi_s,
	z_lo=>q_z_lo_s,
	pc=>q_pc_s,
	mdr=>q_mdr_s, --MDR signal
	inport=>q_inport_s,
	c_sign_extended=>q_c_sign_extended_s,
	s_in=>sel,--select signal
	output=>out_sig); --Bus out
	

phase1_mdr:MDR_unit
	PORT MAP(
		read_sel=>read_sel_s,
		ld =>ld_mdr_s,
		rst_n =>rst_n_s,
		clk =>clk_s,
		BusMuxOut=> q_mdr_s,--:  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		MDataIn=> Mdatain_s,--:  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		Bus_Mux_In=> mdr_s --:  OUT  STD_LOGIC_VECTOR(31 DOWNTO 0));
	);

reg00:reg32bit
	PORT MAP(
	d=>out_sig,
	q=>q00_s,
	ld=>ld00_s,
	rst_n=>rst_n_s,
	clk=>clk_s);

reg01:reg32bit
	PORT MAP(
	d=>out_sig,
	q=>q01_s,
	ld=>ld01_s,
	rst_n=>rst_n_s,
	clk=>clk_s);

reg02:reg32bit
	PORT MAP(
	d=>out_sig,
	q=>q02_s,
	ld=>ld02_s,
	rst_n=>rst_n_s,
	clk=>clk_s);
	
reg03:reg32bit
	PORT MAP(
	d=>out_sig,
	q=>q03_s,
	ld=>ld03_s,
	rst_n=>rst_n_s,
	clk=>clk_s);
	
reg04:reg32bit
	PORT MAP(
	d=>out_sig,
	q=>q04_s,
	ld=>ld04_s,
	rst_n=>rst_n_s,
	clk=>clk_s);

reg05:reg32bit
	PORT MAP(
	d=>out_sig,
	q=>q05_s,
	ld=>ld05_s,
	rst_n=>rst_n_s,
	clk=>clk_s);
	
reg06:reg32bit
	PORT MAP(
	d=>out_sig,
	q=>q06_s,
	ld=>ld06_s,
	rst_n=>rst_n_s,
	clk=>clk_s);
	
reg07:reg32bit
	PORT MAP(
	d=>out_sig,
	q=>q07_s,
	ld=>ld07_s,
	rst_n=>rst_n_s,
	clk=>clk_s);
	
reg08:reg32bit
	PORT MAP(
	d=>out_sig,
	q=>q08_s,
	ld=>ld08_s,
	rst_n=>rst_n_s,
	clk=>clk_s);
	
reg09:reg32bit
	PORT MAP(
	d=>out_sig,
	q=>q09_s,
	ld=>ld09_s,
	rst_n=>rst_n_s,
	clk=>clk_s);
	
reg10:reg32bit
	PORT MAP(
	d=>out_sig,
	q=>q10_s,
	ld=>ld10_s,
	rst_n=>rst_n_s,
	clk=>clk_s);
	
reg11:reg32bit
	PORT MAP(
	d=>out_sig,
	q=>q11_s,
	ld=>ld11_s,
	rst_n=>rst_n_s,
	clk=>clk_s);
	
reg12:reg32bit
	PORT MAP(
	d=>out_sig,
	q=>q12_s,
	ld=>ld12_s,
	rst_n=>rst_n_s,
	clk=>clk_s);
	
reg13:reg32bit
	PORT MAP(
	d=>out_sig,
	q=>q13_s,
	ld=>ld13_s,
	rst_n=>rst_n_s,
	clk=>clk_s);
	
reg14:reg32bit
	PORT MAP(
	d=>out_sig,
	q=>q14_s,
	ld=>ld14_s,
	rst_n=>rst_n_s,
	clk=>clk_s);
	
reg15:reg32bit
	PORT MAP(
	d=>out_sig,
	q=>q15_s,
	ld=>ld15_s,
	rst_n=>rst_n_s,
	clk=>clk_s);

reg_hi:reg32bit
	PORT MAP(
	d=>out_sig,
	q=>q_hi_s,
	ld=>ld_hi_s,
	rst_n=>rst_n_s,
	clk=>clk_s);

reg_lo:reg32bit
	PORT MAP(
	d=>out_sig,
	q=>q_lo_s,
	ld=>ld_lo_s,
	rst_n=>rst_n_s,
	clk=>clk_s);

reg_z_hi:reg32bit
	PORT MAP(
	d=>out_sig,
	q=>q_z_hi_s,
	ld=>ld_z_hi_s,
	rst_n=>rst_n_s,
	clk=>clk_s);	
	
reg_z_lo:reg32bit
	PORT MAP(
	d=>out_sig,
	q=>q_z_lo_s,
	ld=>ld_z_lo_s,
	rst_n=>rst_n_s,
	clk=>clk_s);
	
reg_pc:reg32bit
	PORT MAP(
	d=>out_sig,
	q=>q_pc_s,
	ld=>ld_pc_s,
	rst_n=>rst_n_s,
	clk=>clk_s);
	
reg_inport:reg32bit
	PORT MAP(
	d=>out_sig,
	q=>q_inport_s,
	ld=>ld_inport_s,
	rst_n=>rst_n_s,
	clk=>clk_s);
	
reg_c_sign_extended:reg32bit
	PORT MAP(
	d=>out_sig,
	q=>q_c_sign_extended_s,
	ld=>ld_c_sign_extended_s,
	rst_n=>rst_n_s,
	clk=>clk_s);
END description;
