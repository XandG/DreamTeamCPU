library ieee;
use ieee.std_logic_1164.all;

ENTITY encoder32to5 IS PORT(
    input: IN STD_LOGIC_VECTOR(23 DOWNTO 0);
    sel : OUT STD_LOGIC_VECTOR(4 DOWNTO 0) -- output
);
END encoder32to5;

ARCHITECTURE description OF encoder32to5 IS
BEGIN

process(input)
BEGIN
	case input is
	 when "000000000000000000000001" => sel <="00000";
	 when "000000000000000000000010" => sel <="00001" ;
	 when "000000000000000000000100" => sel <="00010" ;
	 when "000000000000000000001000" => sel <="00011" ;
	 
	 when "000000000000000000010000" => sel <="00100" ;
	 when "000000000000000000100000" => sel <="00101" ;
	 when "000000000000000001000000" => sel <="00110";
	 when "000000000000000010000000" => sel <="00111" ;
	 
	 when "000000000000000100000000" => sel <="01000" ;
	 when "000000000000001000000000" => sel <="01001" ;
	 when "000000000000010000000000" => sel <="01010" ;
	 when "000000000000100000000000" => sel <="01011" ;
	 
	 when "000000000001000000000000" => sel <="01100" ;
	 when "000000000010000000000000" => sel <="01101" ;
	 when "000000000100000000000000" => sel <="01110" ;
	 when "000000001000000000000000" => sel <="01111" ;
	 
	 when "000000010000000000000000" => sel <="10000" ;
	 when "000000100000000000000000" => sel <="10001" ;
	 when "000001000000000000000000" => sel <="10010" ;
	 when "000010000000000000000000" => sel <="10011" ;
	 
	 when "000100000000000000000000" => sel <="10000" ;
	 when "001000000000000000000000" => sel <="10001" ;
	 when "010000000000000000000000" => sel <="10010" ;
	 when "100000000000000000000000" => sel <="10011" ;
	 
	when others => sel<="11111"; -- ERROR SIGNAL
	end case;
	end process;
END description;